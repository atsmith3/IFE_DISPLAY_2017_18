module background(input logic [9:0] disp_x, disp_y,
						output logic [3:0] color,
						output logic draw);
						
	logic [3:0] bg[272][480];
	always_ff begin
		//bg = 
	end
	
	always_comb begin
			draw = 1;
			color = bg[disp_y][disp_x];
	end
	
endmodule