module background
(
    input logic Clk,
    input logic [9:0] DispX, DispY,
    output logic [3:0] color,
    output logic draw
);
logic [3:0] bg[272][480];

always_ff begin
    /*bg = '{'{ , },
            { , }};*/
end

always_comb begin
    draw = 1;
    color = bg[DispX][DispY];
end
endmodule
