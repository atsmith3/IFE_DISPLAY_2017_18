library verilog;
use verilog.vl_types.all;
entity display_tb is
end display_tb;
