module sprite_controller
(
    

);

endmodule
